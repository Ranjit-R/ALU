`define WIDTH 8
`define CMD_WIDTH 4
`define no_of_transactions 10
